module AND_32(out, a, b);
    input [31:0] a, b;
    output[31:0] out;
    
    wire o0, o1, o2, o3, o4, o5, o6, o7, o8, o9, o10, o11, o12, o13, o14, o15;
    wire o16, o17, o18, o19, o20, o21, o22, o23, o24, o25, o26, o27, o28, o29, o30, o31;

    and(o0, a[0], b[0]);
    and(o1, a[1], b[1]);
    and(o2, a[2], b[2]);
    and(o3, a[3], b[3]);
    and(o4, a[4], b[4]);
    and(o5, a[5], b[5]);
    and(o6, a[6], b[6]);
    and(o7, a[7], b[7]);
    and(o8, a[8], b[8]);
    and(o9, a[9], b[9]);
    and(o10, a[10], b[10]);
    and(o11, a[11], b[11]);
    and(o12, a[12], b[12]);
    and(o13, a[13], b[13]);
    and(o14, a[14], b[14]);
    and(o15, a[15], b[15]);
    and(o16, a[16], b[16]);
    and(o17, a[17], b[17]);
    and(o18, a[18], b[18]);
    and(o19, a[19], b[19]);
    and(o20, a[20], b[20]);
    and(o21, a[21], b[21]);
    and(o22, a[22], b[22]);
    and(o23, a[23], b[23]);
    and(o24, a[24], b[24]);
    and(o25, a[25], b[25]);
    and(o26, a[26], b[26]);
    and(o27, a[27], b[27]);
    and(o28, a[28], b[28]);
    and(o29, a[29], b[29]);
    and(o30, a[30], b[30]);
    and(o31, a[31], b[31]);

    assign out[31] = o31;
    assign out[30] = o30;
    assign out[29] = o29;
    assign out[28] = o28;
    assign out[27] = o27;
    assign out[26] = o26;
    assign out[25] = o25;
    assign out[24] = o24;
    assign out[23] = o23;
    assign out[22] = o22;
    assign out[21] = o21;
    assign out[20] = o20;
    assign out[19] = o19;
    assign out[18] = o18;
    assign out[17] = o17;
    assign out[16] = o16;
    assign out[15] = o15;
    assign out[14] = o14;
    assign out[13] = o13;
    assign out[12] = o12;
    assign out[11] = o11;
    assign out[10] = o10;
    assign out[9] = o9;
    assign out[8] = o8;
    assign out[7] = o7;
    assign out[6] = o6;
    assign out[5] = o5;
    assign out[4] = o4;
    assign out[3] = o3;
    assign out[2] = o2;
    assign out[1] = o1;
    assign out[0] = o0;
endmodule
